class tinyalu_env extends uvm_env;
`uvm_component_utils(tinyalu_env)

// Components
tinyalu_agent      agent;
tinyalu_scoreboard scoreboard;
tinyalu_coverage   coverage;

function new(string name, uvm_component parent);
    super.new(name, parent);
endfunction

// Build Phase: Create components
function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    
    agent      = tinyalu_agent::type_id::create("agent", this);
    scoreboard = tinyalu_scoreboard::type_id::create("scoreboard", this);
    coverage   = tinyalu_coverage::type_id::create("coverage", this);
endfunction

// Connect Phase
function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    
    //  Connect Agent -> Scoreboard (Data Checking)
    agent.item_collected_port.connect(scoreboard.item_collected_export);
    
    // Connect Agent -> Coverage (Data Collection)
    agent.item_collected_port.connect(coverage.analysis_export);
endfunction

endclass